module draw_car(
    input clk,
    input resetn,
    input [3:0]COUNTER_X, //Uppercase indicates grid coutner
    input [3:0]COUNTER_Y, //Uppercase indicates grid coutner
    output reg [8:0]colour,
	 output reg draw_done,
    output [7:0]x, //Will go into VGA Input
    output [6:0]y //Will go into VGA Input
    );
    
    wire [8:0]mem_add;
    wire [8:0]colour_car;

    reg [4:0]counter_x;
    reg [4:0]counter_y;
    reg [1:0]one_clk_delay;

    initial begin
        counter_x = 5'b0;
        counter_y = 5'b0;
        one_clk_delay = 1'b0;
        draw_done = 0;
    end

    //Memory Address Translator for 20x20 .mif files
    memory_address_translator_20x20 m1(
                                .x(counter_x), 
                                .y(counter_y), 
                                .mem_address(mem_add) //Connection A
                                ); 

    //.mif-initialized ram with tower image
    ram400x9_car car_unit(
					.address(mem_add), //Connection A
					.clock(clk),
					.data(9'b0),
					.wren(1'b0),
					.q(colour_car)
					);

    always @(posedge clk) begin
        if(!resetn) begin
            counter_x <= 0;
            counter_y <= 0;
            one_clk_delay <= 0;
        end
        else begin
            if(one_clk_delay >= 2'b10)
                one_clk_delay <= 0;
            else
                one_clk_delay <= one_clk_delay + 1;
            
            if(counter_x == 0)
                draw_done <= 0;
                    
            //Loop
            if(one_clk_delay == 2'b10) begin
                counter_x <= counter_x + 1;
                if(counter_x == 5'b10011) begin
                    counter_y <= counter_y + 1;
                    counter_x <= 0;
                end
                    // one_clk_delay <= 0;
            end
        
            //Same as {counter_x, counter_y} >= {19, 19} - i.e. done accessing square memory
            if({counter_x, counter_y} == 10'b1001110011) begin
                draw_done <= 1;
                counter_x <= 0;
                counter_y <= 0;
                one_clk_delay <= 0;
            end
        end
    end

    always @(colour_car) //1 cycle delay from counter_x & counter_y
        colour = colour_car;

    assign x = COUNTER_X * 5'b10100 + counter_x;
    assign y = COUNTER_Y * 5'b10100 + counter_y;
endmodule
